`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date:    Tue Dec  3 14:19:19 2013
// Design Name: 
// Module Name:    netlist_1_EMPTY
//////////////////////////////////////////////////////////////////////////////////
module netlist_1_EMPTY(DIP, LED, LCDDATA, CLK, CLK_33MHZ_FPGA, nRST, BTN_N, BTN_E, BTN_S, BTN_W, BTN_C, LED_N, LED_E, LED_S, LED_W, LED_C, RS, RW, EN);
  input [7:0] DIP;
  output [7:0] LED;
  inout  [3:0] LCDDATA;
  input CLK;
  input CLK_33MHZ_FPGA;
  input nRST;
  input BTN_N;
  input BTN_E;
  input BTN_S;
  input BTN_W;
  input BTN_C;
  output LED_N;
  output LED_E;
  output LED_S;
  output LED_W;
  output LED_C;
  output RS;
  output RW;
  output EN;


endmodule
